module archive_00001(a, b, y);
input [4+5+6+4+5+6-1:0] a;
wire [3:0] a0 = a[4-1:0];
wire [4:0] a1 = a[4+5-1:4];
wire [5:0] a2 = a[4+5+6-1:4+5];
wire signed [3:0] a3 = a[4+5+6+4-1:4+5+6];
wire signed [4:0] a4 = a[4+5+6+4+5-1:4+5+6+4];
wire signed [5:0] a5 = a[4+5+6+4+5+6-1:4+5+6+4+5];
input [4+5+6+4+5+6-1:0] b;
wire [3:0] b0 = b[4-1:0];
wire [4:0] b1 = b[4+5-1:4];
wire [5:0] b2 = b[4+5+6-1:4+5];
wire signed [3:0] b3 = b[4+5+6+4-1:4+5+6];
wire signed [4:0] b4 = b[4+5+6+4+5-1:4+5+6+4];
wire signed [5:0] b5 = b[4+5+6+4+5+6-1:4+5+6+4+5];
output [4+5+6+4+5+6-1:0] y;
wire [3:0] y0;
wire [4:0] y1;
wire [5:0] y2;
wire signed [3:0] y3;
wire signed [4:0] y4;
wire signed [5:0] y5;
assign y = {y0,y1,y2,y3,y4,y5};
assign y0 = ((^(^((a5)))));
assign y1 = ((((((a3))))));
assign y2 = {((({a5,b4,b2}*(b0^b3)))),({((a4)*(b5))}),{({b0,a0}&&{(a4^a3)})}};
assign y3 = ({(({(b1||b0)})^~((a5^b3)&&(a0)))}<<{{a4,a2,a2},(a1^a2),{b3,a3,b0}});
assign y4 = (~^{a3,b2});
assign y5 = (+((~^(~((-(|a2))&(a3*b0))))^~(((b4|a3)*(a2>>>a1))>>>((a4>>a2)^(~b5)))));
endmodule
